library IEEE; 
use IEEE.STD_LOGIC_1164.all; 

package projectPackage is
    type FEATURE_type is array (integer range <>) of std_logic_vector(31 downto 0);
    type CENTROID_type is array (integer range <>) of std_logic_vector(31 downto 0);

end projectPackage; 

package body projectPackage is 

end projectPackage; 